//                              -*- Mode: Verilog -*-
// Filename        : adxl362_accelerometer.v
// Description     : ADXL362 Accelerometer Module
// Author          : Philip Tracton
// Created On      : Thu Jun 23 20:53:26 2016
// Last Modified By: Philip Tracton
// Last Modified On: Thu Jun 23 20:53:26 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!

module adxl362_accelerometer (/*AUTOARG*/ ) ;
   
endmodule // adxl362_accelerometer
