//                              -*- Mode: Verilog -*-
// Filename        : adxl362_fifo.v
// Description     : ADXL362 512 element FIFO
// Author          : Philip Tracton
// Created On      : Thu Jun 23 20:54:03 2016
// Last Modified By: Philip Tracton
// Last Modified On: Thu Jun 23 20:54:03 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!

module adxl362_fifo (/*AUTOARG*/ ) ;
   
endmodule // adxl362_fifo
