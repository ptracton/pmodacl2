//                              -*- Mode: Verilog -*-
// Filename        : spi_tasks.v
// Description     : SPI Tasks
// Author          : Philip Tracton
// Created On      : Fri Jul  8 21:12:20 2016
// Last Modified By: Philip Tracton
// Last Modified On: Fri Jul  8 21:12:20 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!

module spi_tasks (/*AUTOARG*/ ) ;
   
endmodule // spi_tasks
