//                              -*- Mode: Verilog -*-
// Filename        : adxl362_testbench.v
// Description     : Testbench for proving ADXL362 Model works
// Author          : Philip Tracton
// Created On      : Wed Jun 22 21:42:09 2016
// Last Modified By: Philip Tracton
// Last Modified On: Wed Jun 22 21:42:09 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!

module adxl362_testbench (/*AUTOARG*/ ) ;


   
   
endmodule // adxl362_testbench
