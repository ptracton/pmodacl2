//                              -*- Mode: Verilog -*-
// Filename        : adxl362_temperature.v
// Description     : ADXL362 Temperature Sensor
// Author          : Philip Tracton
// Created On      : Thu Jun 23 20:55:46 2016
// Last Modified By: Philip Tracton
// Last Modified On: Thu Jun 23 20:55:46 2016
// Update Count    : 0
// Status          : Unknown, Use with caution!

module adxl362_temperature (/*AUTOARG*/ ) ;
   
endmodule // adxl362_temperature
